module testbench

endmodule
